module armreduced(
	input clk,
	input reset,
	output[31:0] pc,
	input[31:0] inst,
	input nIRQ,
	output[3:0] be,
	output[31:0] memaddr,
	output memwrite,
	output memread,
	output[31:0] writedata,
	input[31:0] readdata
	);
	assign be = 4'b1111; // default
	assign memread = 'b1; // default
	
	RegisterFile registerfile();
	ALU alu();
	ControlUnit controlunit();
	Extend extend();
	
	always@(posedge clk or negedge reset) begin
		
	end
	
endmodule
