module RegisterFile(
	);
	
	reg[31:0] register[15:0]; 	

endmodule
